    Mac OS X            	   2  �     �                                    ATTRQt�  �   �  �                  �   C  com.apple.quarantine     b  %com.apple.metadata:kMDItemWhereFroms 0001;5886cefd;Google\x20Chrome;6A5DADF9-79C4-443B-A51B-FCF1D0BD22EBbplist00�_�https://connect.ubc.ca/bbcswebdav/pid-3824145-dt-content-rid-18667172_1/courses/SIS.UBC.CPEN.391.201.2016W2.74350/SIS.UBC.CPEN.391.201.2016W2.74350_ImportedContent_20161011050002/ACIA_Clock.vhd_jhttps://connect.ubc.ca/webapps/blackboard/content/listContent.jsp?course_id=_87470_1&content_id=_3824082_1   �                           <                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                  This resource fork intentionally left blank                                                                                                                                                                                                                            ��