    Mac OS X            	   2  �     �                                    ATTR3zA  �   �  �                  �   C  com.apple.quarantine     _  %com.apple.metadata:kMDItemWhereFroms 0001;5886cf00;Google\x20Chrome;FDE2F1B1-9623-409F-8C6E-E435187660EDbplist00�_�https://connect.ubc.ca/bbcswebdav/pid-3824145-dt-content-rid-18667174_1/courses/SIS.UBC.CPEN.391.201.2016W2.74350/SIS.UBC.CPEN.391.201.2016W2.74350_ImportedContent_20161011050002/ACIA_TX.vhd_jhttps://connect.ubc.ca/webapps/blackboard/content/listContent.jsp?course_id=_87470_1&content_id=_3824082_1   �                           9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     This resource fork intentionally left blank                                                                                                                                                                                                                            ��