    Mac OS X            	   2  �     �                                    ATTR���  �   �  �                  �   C  com.apple.quarantine     a  %com.apple.metadata:kMDItemWhereFroms 0001;5886cefc;Google\x20Chrome;302C2969-E4BC-44C4-B3EA-59153A018AB0bplist00�_�https://connect.ubc.ca/bbcswebdav/pid-3824145-dt-content-rid-18667171_1/courses/SIS.UBC.CPEN.391.201.2016W2.74350/SIS.UBC.CPEN.391.201.2016W2.74350_ImportedContent_20161011050002/ACIA_6850.vhd_jhttps://connect.ubc.ca/webapps/blackboard/content/listContent.jsp?course_id=_87470_1&content_id=_3824082_1   �                           ;                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                   This resource fork intentionally left blank                                                                                                                                                                                                                            ��