    Mac OS X            	   2  �     �                                    ATTRK��  �   �  �                  �   C  com.apple.quarantine     d  %com.apple.metadata:kMDItemWhereFroms 0001;5886cf03;Google\x20Chrome;0D112683-F0CA-4003-B9A9-92E5D7A52ED4bplist00�_�https://connect.ubc.ca/bbcswebdav/pid-3824145-dt-content-rid-18673211_1/courses/SIS.UBC.CPEN.391.201.2016W2.74350/SIS.UBC.CPEN.391.201.2016W2.74350_ImportedContent_20161011050002/Register3Bit.vhd_jhttps://connect.ubc.ca/webapps/blackboard/content/listContent.jsp?course_id=_87470_1&content_id=_3824082_1   �                           >                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                This resource fork intentionally left blank                                                                                                                                                                                                                            ��