    Mac OS X            	   2  �     �                                    ATTR~�WL  �   �  �                  �   C  com.apple.quarantine     _  %com.apple.metadata:kMDItemWhereFroms 0001;5886ceff;Google\x20Chrome;B48CC98F-E993-4657-BB9D-6D57429EC903bplist00�_�https://connect.ubc.ca/bbcswebdav/pid-3824145-dt-content-rid-18667173_1/courses/SIS.UBC.CPEN.391.201.2016W2.74350/SIS.UBC.CPEN.391.201.2016W2.74350_ImportedContent_20161011050002/ACIA_RX.vhd_jhttps://connect.ubc.ca/webapps/blackboard/content/listContent.jsp?course_id=_87470_1&content_id=_3824082_1   �                           9                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                     This resource fork intentionally left blank                                                                                                                                                                                                                            ��