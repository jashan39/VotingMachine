    Mac OS X            	   2  �     �                                    ATTR
�%  �   �   C                  �   C  com.apple.quarantine 0001;5886cf46;Google\x20Chrome;76D73BB4-F23F-41E6-95B1-211CAF102BF7                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                    This resource fork intentionally left blank                                                                                                                                                                                                                            ��